    .INIT_00(256'h0000001dcff1f0000000000bc1b0b01d00000034a3a1f0000000001dcff0b01c),
    .INIT_01(256'h00000034a3a0b0020000001dcff2023b0000000bc1a2023200000034a3436017),
    .INIT_02(256'h0000000bc1c0b00200000034a34202440000001dcff323770000000bc1d1d002),
    .INIT_03(256'h0000000bd202b40f000000250002024d00000034a3a323770000001dcff1d003),
    .INIT_04(256'h00000020a34010400000000bc172b04f00000032a182b08f0000001dd002b20f),
    .INIT_05(256'h00000020a46010080000000bc202d01000000020a40010200000000bc162d010),
    .INIT_06(256'h0000000bc192b80f00000032a212d0100000001dd00010040000000bd212d010),
    .INIT_07(256'h0000000bc210101000000020a402d0100000000bc180108000000020a342b10f),
    .INIT_08(256'h00000032a2a1d0010000001dd000b0320000000bd2220b0800000020a462d010),
    .INIT_09(256'h00000020a402f01e0000000bc1a0100100000020a34220080000000bc1b326c5),
    .INIT_0A(256'h0000001dd0011d010000000bd230bf1200000020a460be110000000bc220bd10),
    .INIT_0B(256'h0000000bc1c2fe1100000020a342fd100000000bc1d13f0000000032a3313e00),
    .INIT_0C(256'h000000250000b00f00000020a4620e7a0000000bc232ff1200000020a4003f03),
    .INIT_0D(256'h0000002086b030fc000000208930b03b000000208b72f00f000000208dd03007),
    .INIT_0E(256'h000000208d73646d000000208b31c0e00000002500003efc000000208930be0e),
    .INIT_0F(256'h000000250001d00100000020891324450000002086b1d000000000208930b001),
    .INIT_10(256'h0000002086b1d003000000208933244d000000208d71d002000000208b332449),
    .INIT_11(256'h000000208db20be5000000208c720a7a0000002500020b910000002089332451),
    .INIT_12(256'h0000002500020be50000002089120a810000002086b20b940000002089322454),
    .INIT_13(256'h0000002b08e20be50000002b1bb20a8b0000002b21a20b970000002bec922454),
    .INIT_14(256'h00000001c0020be50000002500020a970000002005c20b9a00000020bd122454),
    .INIT_15(256'h00000020a651f00000000001c100b017000000250001d00000000020a650b016),
    .INIT_16(256'h000000250001f00000000020a650b01900000001c071f000000000250000b018),
    .INIT_17(256'h00000001c011f000000000250000b01b00000020a651f00000000001c0d0b01a),
    .INIT_18(256'h00000020a651f00000000001c040b01d000000250001f00000000020a650b01c),
    .INIT_19(256'h00000001f002093000000001e002091100000001d002246d0000002500036466),
    .INIT_1A(256'h00000020b60209020000000110001004000000010802094100000020b6920891),
    .INIT_1B(256'h0000002b00a0b0020000002b3892023b000000250002023200000020a7422008),
    .INIT_1C(256'h000000250000b00200000020bd1202440000002b08e324770000002b63b1d002),
    .INIT_1D(256'h0000002b08e2b40f0000002b37b2024d0000002b00a324770000002b2091d003),
    .INIT_1E(256'h0000002b6490104000000020a622b04f000000250002b08f00000020bd12b20f),
    .INIT_1F(256'h00000020bd1010080000002b08e2d0100000002b5bb010200000002b62a2d010),
    .INIT_20(256'h00000020a4c2b80f00000020b022d01000000020a4c01004000000250002d010),
    .INIT_21(256'h0000002b5bb010100000002b62a2d0100000002b6490108000000020a622b10f),
    .INIT_22(256'h00000020a4c2b10f000000250002b80f00000020bd120b080000002b08e2d010),
    .INIT_23(256'h00000020a4c2d01000000020b020101000000020a4c2d01000000020b0201080),
    .INIT_24(256'h0000002b5bb220080000002b62a209300000002b6492090200000020a6201002),
    .INIT_25(256'h00000020a4c0d004000000250000900e00000020bd12f0320000002b08e01000),
    .INIT_26(256'h00000020a4c0901800000020b022f00700000020a4c0901700000020b02324c3),
    .INIT_27(256'h0000002b6490901a00000020a622f00900000020a4c0901900000020b022f008),
    .INIT_28(256'h00000020bd1090160000002b08e2f00b0000002b5bb0901b0000002b62a2f00a),
    .INIT_29(256'h0000002b10a1d00a0000002b6490300f00000020a5f2b04e000000250002f033),
    .INIT_2A(256'h0000002b6c93261b00000020bd10d0020000002b08e090020000002bdfb364ad),
    .INIT_2B(256'h00000020bd12261b0000002b08e364b00000002bebb1d00e0000002b10a2261c),
    .INIT_2C(256'h00000020b8503c0f00000001ccc0bc0700000020a4c364ba000000250001d00b),
    .INIT_2D(256'h0000002b6492086b00000020a5f2089300000020a4c208d300000020af62dc01),
    .INIT_2E(256'h00000020bd1364be0000002b08e1d00f0000002bdfb220030000002b10a20891),
    .INIT_2F(256'h0000002b08e326420000002bebb1d00c0000002b10a2262d0000002b6c9208b7),
    .INIT_30(256'h00000001cd80900d00000020a4c22619000000250003264200000020bd10d008),
    .INIT_31(256'h00000001ccc1d04f00000020a4c0900600000020af63661b00000020b850d020),
    .INIT_32(256'h00000020a5f3261b00000020a4c0d00200000020af60900200000020b85364cd),
    .INIT_33(256'h0000002b08e208d50000002bdfb364d90000002b10a1d0530000002b6492261c),
    .INIT_34(256'h0000002bebb209390000002b10a013000000002b6c90b20200000020bd120891),
    .INIT_35(256'h00000020a4c364d3000000250001c32000000020bd1113010000002b08e20948),
    .INIT_36(256'h00000020a4c208d300000020af6364f000000020b851d05200000001ce42261a),
    .INIT_37(256'h00000020a4c3661900000020af61d02000000020b850900600000001cd8208e8),
    .INIT_38(256'h00000020a4c1d03000000020af60900600000020b85208e800000001ccc20893),
    .INIT_39(256'h0000002bdfb090060000002b10a208e80000002b6492089d00000020a5f36619),
    .INIT_3A(256'h0000002b10a001000000002b6c92d00100000020bd13a6190000002b08e2085e),
    .INIT_3B(256'h000000250002200300000020bd1208910000002b08e208e50000002bebb2087c),
    .INIT_3C(256'h0000002b08e2262d0000002b47b208b70000002b22a364f40000002b1c91d044),
    .INIT_3D(256'h0000002b22a208e80000002b489208cb000000250003651b00000020bd11d04e),
    .INIT_3E(256'h000000250002089300000020bd1366190000002b08e1d0200000002b57b09006),
    .INIT_3F(256'h0000002b08e2fa080000002b6bb3a6190000002b66a208810000002b5c90120a),
    .INIT_40(256'h0000002b66a2fe330000002b6c92fd0b000000250002fc0a00000020bd12fb09),
    .INIT_41(256'h0000002500014a0600000020bd13a6190000002b08e208810000002b7bb01201),
    .INIT_42(256'h000000010800bb0800000020a4c14a0600000020b0214a0600000020a4c14a06),
    .INIT_43(256'h000000250000bf3300000020a6e0be0b00000020b600bd0a000000011010bc09),
    .INIT_44(256'h00000020af62085700000020b852085700000001c0e2085700000020a4c20857),
    .INIT_45(256'h00000020a4c2fd0a000000250002fc0900000020a532fb0800000020a4c2fa07),
    .INIT_46(256'h00000020a4c1d05400000020af62265300000020b852ff3300000001c1e2fe0b),
    .INIT_47(256'h00000020af60900600000020b85208e800000001c0e208d700000020a5336588),
    .INIT_48(256'h00000020a4c0120a000000250002089300000020a533661900000020a4c1d020),
    .INIT_49(256'h00000020a4c2fb0900000020af62fa0800000020b853a61900000001c2e20881),
    .INIT_4A(256'h00000020af60120100000020b852fe3300000001c1e2fd0b00000020a532fc0a),
    .INIT_4B(256'h00000020b8514a0600000001c0e3a61900000020a533a61900000020a4c20881),
    .INIT_4C(256'h000000250002fa0700000020a5314a0600000020a4c14a0600000020af614a06),
    .INIT_4D(256'h0000001d0030bd0a00000032b3b0bc090000001d0020bb080000000b0020ba07),
    .INIT_4E(256'h00000020b102085700000032b3f208570000001d0040bf3300000032b3d0be0b),
    .INIT_4F(256'h00000020b232fb0800000022b402fa0700000020b172085700000022b4020857),
    .INIT_50(256'h00000001c0e2ff3300000020a4c2fe0b000000250002fd0a0000000b0022fc09),
    .INIT_51(256'h000000250003256a00000020a4c1df0c00000020af62fb3f00000020b852fa3e),
    .INIT_52(256'h00000020af60ba3300000020b852261900000001c1a3254b00000020a4c0df08),
    .INIT_53(256'h00000020af62085000000020b852085000000001c0e2085000000020a4c2fa13),
    .INIT_54(256'h00000001c262fe0e00000020a4c2fd0d000000250002fc0c00000020a4c20850),
    .INIT_55(256'h00000001c1a0bd1000000020a4c2089100000020af620d8500000020b852ff0f),
    .INIT_56(256'h00000001c0e2089d00000020a4c208b500000020af60bf1200000020b850be11),
    .INIT_57(256'h000000250002086b00000020a4c00ce000000020af62086b00000020b8500cf0),
    .INIT_58(256'h0000002d108208720000002d0080bc3f0000002b4192086b0000002b00a00cd0),
    .INIT_59(256'h0000002d1080bc3e0000002d008208e50000002b2592087c0000002b00a20872),
    .INIT_5A(256'h0000002dc08208500000002b289208500000002b00a22619000000250002086b),
    .INIT_5B(256'h0000002500003e030000002df08208500000002de08208500000002dd082fe13),
    .INIT_5C(256'h00000009d0820e7a00000009c082fe120000002b2892fd110000002b00a2fc10),
    .INIT_5D(256'h0000002d10a0bd0e000000250000be0d00000009f080bf0c00000009e0820891),
    .INIT_5E(256'h0000002de082086b0000002dd0800cd00000002dc082086b0000002d0090bc0f),
    .INIT_5F(256'h0000002d0092086b0000002d10a00cf0000000250002086b0000002df0800ce0),
    .INIT_60(256'h00000009f082087c00000009e082087200000009d082087200000009c080bc3f),
    .INIT_61(256'h0000002d10a22619000000011022086b000000010500bc3e00000025000208e5),
    .INIT_62(256'h00000020a6e0d00400000025000090020000002dc08365a60000002d0091d058),
    .INIT_63(256'h00000020a740900600000020b69208e800000025000208df00000020b703e5a6),
    .INIT_64(256'h000000250000120800000020b9d2089300000020a4c36619000000250001d020),
    .INIT_65(256'h00000020b482fa34000000250002089100000020b9d3a61900000020b4220881),
    .INIT_66(256'h00000020b9d0bc3400000020b522fd3b000000250002fc3600000020b9d2fb35),
    .INIT_67(256'h00000020b6001a01000000011000bf3b000000010200be36000000250000bd35),
    .INIT_68(256'h0000000bc0c09c070000000bd0d208080000000be0e208280000000bf0f01b00),
    .INIT_69(256'h000000010803661b00000020b911d051000000250002261900000020b8e2086b),
    .INIT_6A(256'h000000011001d020000000010000900600000020b60208e800000001101208d1),
    .INIT_6B(256'h000000250002088100000020aa50120a00000020b8e2089300000020b7e36619),
    .INIT_6C(256'h000000011012fc0a000000010802fb0900000020b422fa0800000020b943a619),
    .INIT_6D(256'h00000020b7e208810000000110001201000000010042fe3300000020b602fd0b),
    .INIT_6E(256'h00000020b9714a060000002500014a0600000020ab114a0600000020b8e3a619),
    .INIT_6F(256'h00000020b600bd0a000000011010bc09000000010800bb0800000020b4814a06),
    .INIT_70(256'h00000020b8e2085700000020b7e20857000000011000bf33000000010080be0b),
    .INIT_71(256'h00000020b522fb0800000020b9a2fa07000000250002085700000020ac220857),
    .INIT_72(256'h0000000100c2ff3300000020b602fe0b000000011012fd0a000000010802fc09),
    .INIT_73(256'h00000020ad7325d100000020b8e0df0800000020b7e325db000000011001df0c),
    .INIT_74(256'h00000036bd1208500000000d008208500000000900e2ff130000002500022619),
    .INIT_75(256'h00000032bd52fd0d0000000d0022fc0c0000000900e208500000002500020850),
    .INIT_76(256'h00000032bd9208500000000d002225f00000000900f2ff0f000000250002fe0e),
    .INIT_77(256'h00000032bdd208500000000d00220850000000090102fe130000002500020850),
    .INIT_78(256'h00000032be12fe120000000d0022fd11000000090112fc100000002500003e03),
    .INIT_79(256'h0000002f11618c00000000011000b206000000370010b105000000250000b004),
    .INIT_7A(256'h0000002f11a20e7a0000002f1193e6190000002f1181ae200000002f1171ad10),
    .INIT_7B(256'h000000010a2225f00000002f11d2f40f0000002f11c034070000002f11b0b40f),
    .INIT_7C(256'h00000011001325fa0000002b00b1d0000000002b00a0b0130000002b6c920b34),
    .INIT_7D(256'h0000001d0ff3260000000020c5a1d00200000020c00325fd00000020bfb1d001),
    .INIT_7E(256'h00000009c0820a7a0000002500020b91000000370003260500000036bf31d003),
    .INIT_7F(256'h000000250002260500000009f0820a8100000009e0820b9400000009d0822605),
    .INITP_00(256'h38023bba2aa53b0d1d341732aaaaa6a51132b28d28a597a3ba15a1be98bbbd12),
    .INITP_01(256'h243fada0003236372c21a40db1853e95b43ea92a3b1e06ac15afb035323d8385),
    .INITP_02(256'ha8be00a0b48f2fb800a7a708a92f1005bc90b525af2b2eb8861621ababa38a3a),
    .INITP_03(256'h9fbc289c3704aa80ba229a29b31e24951e30bd11bd9086342b010fa900a7b48a),
    .INITP_04(256'h229804868701008a1b211b23b399209c830d830807b708bc2b9cb0029b1b9aaf),
    .INITP_05(256'h2c15a105083335ac289480b2312c0aa687b79021979cb33aaba89d3007273f84),
    .INITP_06(256'h0424ada880a62baa0fbc0eb61dbd138abcb4ada30a18a925af0aa4b021863f1e),
    .INITP_07(256'hbebc3995a7803eb7b889ae003c193f26208abf1e210b01313320af1b882f2523),
    .INITP_08(256'h2f25361f8f2aa6a688af1206af2dba8a2e8f369004900890bc01b88bb289a98b),
    .INITP_09(256'h110c8a80170b9f118b1d95352a0e90b537b51b87b4aba51b0fa422a890a79a01),
    .INITP_0A(256'h249d2db3bf022ea7320ea624bf08aa0a2fad3a09a5212687b1172a263108a4b3),
    .INITP_0B(256'h89372482342590022e249c373d98060f3515363d920c0724bb1b9a84bd1bb31f),
    .INITP_0C(256'hbd0f3c2325af2b293c2221be392f042d16b82d399fa0978fa59915ac1b3cbb1d),
    .INITP_0D(256'h369004af32bc893ebe9b39b69584b8a6ab0b303d0b233f150aafaab3be9f13a1),
    .INITP_0E(256'h0cbb1b2610bd802193371326a4bd92aa333ca81da9b598082b3fa63231b308bf),
    .INITP_0F(256'ha29331309121b7a79e96b9950010148c0399921d96858a8a071d27b003b10935),
