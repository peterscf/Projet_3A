    .INIT_00(256'h022dfd208f620a4c011f010504025000013a00208f020b8e01390020b0803cff),
    .INIT_01(256'h032e0d22008201fc01cf50209300110000b2382090201010001f0001000201f8),
    .INIT_02(256'h011f012500025000013a003680820b770139000d080010140108200900d01100),
    .INIT_03(256'h032e15250000110001cf303680c01014001f000d040201f8022e060900d20b42),
    .INIT_04(256'h011f010b21520b7701380001300010140139000150a0110001180101440201fc),
    .INIT_05(256'h003a03143000101802f91114200201f802f8100d01020b48022e0e0b01425000),
    .INIT_06(256'h004a000300701018014006143000110001400614200201fc00b0130d00801100),
    .INIT_07(256'h00bd3014106201f80250003a82120b52037000190012500002fa120110120b77),
    .INIT_08(256'h0019002d30a0101c00180012350201fc00b237102400110000be312281d0101c),
    .INIT_09(256'h032e2d2500020b7e01cf200201025000001f000900820b77001a002d20901100),
    .INIT_0A(256'h011f012de0703cff013a002080c03dfe0129e02df0703eff0108d02080c03fff),
    .INIT_0B(256'h01df002dc0705c00003ff02080c05d0100bf392dd0705e00022e262080c05f00),
    .INIT_0C(256'h01df022da07201f800b23c2080c20a4c001f002db0725000032e3a2080c20b8e),
    .INIT_0D(256'h013a00013000110001390001500202270108200146c01100032e3a2500001010),
    .INIT_0E(256'h00b2381420020b42001f000d01025000022e330b01420b77011f010b21501014),
    .INIT_0F(256'h0108201430020227032e44142000110001cf000d0080101400b03714300201f8),
    .INIT_10(256'h022e3c3a84625000011f011900120b77013a0001101010140139000300701100),
    .INIT_11(256'h032e4d123500110001cf50102400101800b20322842201f8001f001410620b48),
    .INIT_12(256'h011f010601020b77013a0009008010180139002d209011000108202d30a20227),
    .INIT_13(256'h032e55250000101c01cf302d008201f8001f002d20920b52022e462d30a25000),
    .INIT_14(256'h011f0114d000110001380014c000101c01390014b002022701180114a0601100),
    .INIT_15(256'h003a0314f0e2f03202f911250000100002f81014f0025000022e4e14e0020b77),
    .INIT_16(256'h004a0014b083228901400614c080d00801400614d080901100b01314e082f01e),
    .INIT_17(256'h020e73390001d004025000110b932265037000250001d00802fa1214a0809012),
    .INIT_18(256'h0096083e8681d001009508190113227702f503390001d002009508190e93226e),
    .INIT_19(256'h009608250000900f009508190f62f00102f605390000100002f5041100732280),
    .INIT_1A(256'h00960820872362e300950800c000d02002f63125000362e302f5301100a0d040),
    .INIT_1B(256'h0096082087c2f001009508208720100102f638208e5362cd02f5372087c0d080),
    .INIT_1C(256'h0015ef14c060d00402500001100362e302f606250000d00802f53c208e50900f),
    .INIT_1D(256'h02d60a14c060100202d50914100362cd00110014c060d01000160714100362e3),
    .INIT_1E(256'h020e5f25000362e3037001141000d04002500014c060901002d10b141002f001),
    .INIT_1F(256'h02f83411130362cd00ba12111070d08000b9113a87f362e300b8101d10a0d020),
    .INIT_20(256'h00bd37090060d008001200208e80901002fa3601a002f00102f9352500001003),
    .INIT_21(256'h01a940208500d01001883001104362e300b431390000d00400b3302085e362e3),
    .INIT_22(256'h02f83400100362c901120104a000d08003ae91368870900e01ba0019101362cd),
    .INIT_23(256'h032ebd36882362c301c2d0192010d02002fa36208e5362c602f9352087c0d040),
    .INIT_24(256'h00ba36011200d00400b935228e50900e00b8340110d362c0022e86250000d010),
    .INIT_25(256'h0094080113e2b04e001300228e52f0330012000115f0901602f20f228e53229c),
    .INIT_26(256'h01b90001133222af018840228e5362ae032f4f011311d00e01d401228e50300f),
    .INIT_27(256'h0133000113109006011201228e5362ae03aea4011300d02001ba00228e50900d),
    .INIT_28(256'h022e97011331d05302fa36228e5222af02f93501132362a302f834228e51d049),
    .INIT_29(256'h02f30e011350b20200ba36228e52089100b93501134208d500b834228e5362ae),
    .INIT_2A(256'h00b50d011371c32000b40c228e51130102f80c011362093902f20d228e501300),
    .INIT_2B(256'h01460801139208c100b30e228e52200800b70f011382093000b60e228e5362a9),
    .INIT_2C(256'h014700011420b002014308228e52020c0147000114120203014608228e520891),
    .INIT_2D(256'h014006011440b002014006228e52021500b01301143322bb02f70e228e51d002),
    .INIT_2E(256'h0370000114620b0802f00f228e52021e01400601145322bb014006228e51d003),
    .INIT_2F(256'h01d40001148220080034f0228e52093000b4390114720902025000228e501000),
    .INIT_30(256'h0188400114a2b20e001200228e5222e100b43c0114901080032ef3228e52b10e),
    .INIT_31(256'h0112010114c0102003aece228e52b40e01ba000114b222e101b900228e501040),
    .INIT_32(256'h01d2020114e0101002fa36228e52b80e02f9350114d20b3402f834228e5222e1),
    .INIT_33(256'h00b935011501d00000b834228e50b001022ec30114f20b34032ef3228e5222e1),
    .INIT_34(256'h019402011521d00200b43c228e5322d902f20f011511d00100ba36228e5322d7),
    .INIT_35(256'h03ef4f011542b80f01ba00228e5322de01b900011531d003018840228e5322db),
    .INIT_36(256'h00b20f011560108000ba36228e5222e000b935011552b10f00b834228e5222e0),
    .INIT_37(256'h014808011582d01001490e228e50101000330101157222e0000380228e52d010),
    .INIT_38(256'h0149080115a20203000390228e5223e202f80d011592f01e02f30c228e501008),
    .INIT_39(256'h01420625000322ed0143082d1061d002014200208ec0b002014908228e52020c),
    .INIT_3A(256'h01400625000322ed00b013368e81d0030013020d0200b00202f20e0900d20215),
    .INIT_3B(256'h00430025000322f6014006368ec1d0000140060d0100b0010140060900d2021e),
    .INIT_3C(256'h00b43809000322fc025000250001d00203700003060322f902f30f090001d001),
    .INIT_3D(256'h01ba00031602b20f01b900001002b40f01884025000323010012000309f1d003),
    .INIT_3E(256'h02f935208bb2230502f8342d1002b04f011201041002b08f03af00208f322305),
    .INIT_3F(256'h022ef52086a2d010032f22208f00102001c2d0208932d01002fa36208b501040),
    .INIT_40(256'h02f20f0319f0100400ba36001002d01000b935250000100800b8342089122305),
    .INIT_41(256'h01b900208d50982f0188402d1002f01e019402041000100100b438208f02d010),
    .INIT_42(256'h00b9351d0011d00000b8340b0320b00103ef4f208930b23701ba00208b519801),
    .INIT_43(256'h02f30c208911d0020013002086a3231e00b20f208f31d00100ba363292c32313),
    .INIT_44(256'h01490820893010a0014908208b53233c000390208d51d00302f80d250003232c),
    .INIT_45(256'h02f20e2500003f070142002089120b8b0143082086a20b600142000100201102),
    .INIT_46(256'h014006041002ff0f014006208f02fe0e00b0130319f2fd0d001303001002fc0c),
    .INIT_47(256'h02f30f2091820b020043000100020a4c014006250002234e0140062d10020b91),
    .INIT_48(256'h001200208b520b6000b403208d5011020250002d103010a00370000b13220a4c),
    .INIT_49(256'h03af2d3292c2fd0d01ba001d0012fc0c01b9000b03203f070188402089320b8b),
    .INIT_4A(256'h02fa36250002235102f9352089120b9402f8342086a2ff0f011201010402fe0e),
    .INIT_4B(256'h00ba362500020b0200b9352089120a4c00b8342086a20b02022f240102020a4c),
    .INIT_4C(256'h018840208cd20b60019402329370110200b4031d000010a002f20f208f320a4c),
    .INIT_4D(256'h00b834208c12fd0d03ef4f250002fc0c01ba002089303f0701b9002089720b8b),
    .INIT_4E(256'h001300208932235400b20f208cb20b9700ba36208d52ff0f00b935229342fe0e),
    .INIT_4F(256'h0149082090720b020003902089120a4c02f80d2086b20b0202f30c00c3020a4c),
    .INIT_50(256'h01420020893010a0014308208c120a4c014200208d320b02014908208fb20a4c),
    .INIT_51(256'h0140062500003f0700b0132089120b8b0013042086b20b6002f20e0bc3a01102),
    .INIT_52(256'h0043002089d2ff0f014006208932fe0e014006208bb2fd0d014006208c92fc0c),
    .INIT_53(256'h0012ff0bc0520be50250002086b20a7a0370000bc062235702f30f2089d20b9a),
    .INIT_54(256'h02f20f208912235902f20e2086b20be502f20d0bc0420a8102f20c2086b22359),
    .INIT_55(256'h00b0162089320a97001300208b322359025000208d720be50370002099e20a8b),
    .INIT_56(256'h02f117209b00b01702f0163a95d1d000020f730d5040b01600b1170950220be5),
    .INIT_57(256'h00b11909e1e0b01900b01809d1d1f00000130109c1c0b01802f220229741f000),
    .INIT_58(256'h02f22114b060b01b02f11914b061f00002f0180bb130b01a020f7309f1f1f000),
    .INIT_59(256'h020f7313f000b01d00b11b13e001f00000b01a13d000b01c00130210cb01f000),
    .INIT_5A(256'h0013032fc341100102f2222fd350b03a02f11b2fe363638e02f01a2ff3b1f000),
    .INIT_5B(256'h02f01c2086b0b002020f730bc362023b00b11d2086b2023200b01c0bc3b2f03a),
    .INIT_5C(256'h0012002086b0b0020250000bc342024402f2232086b3237702f11d0bc351d002),
    .INIT_5D(256'h014006208932b40f031000208b32024d01f1ff208b53237701d0ff208911d003),
    .INIT_5E(256'h0141002299201040014006209b02b04f0140063a97c2b08f0140060d5042b20f),
    .INIT_5F(256'h01400e0bf3b0100801400e0be362d0100141000bd35010200140060bc342d010),
    .INIT_60(256'h025000208082b80f00b224208282d01001003001b000100401400e01a042d010),
    .INIT_61(256'h022ffd2080801010022ffd09e072d010022ffd2080801080022ffd09f072b10f),
    .INIT_62(256'h022ffd2086b1d001022ffd09c070b032022ffd2080820b08022ffd09d072d010),
    .INIT_63(256'h022ffd2086b323dd022ffd00ce01d800022ffd2086b22008022ffd00cd0326c5),
    .INIT_64(256'h022ffd208b52f035022ffd208910b017022ffd2086b2f034022ffd00cf00b016),
    .INIT_65(256'h022ffd01c002f03b022ffd2089d0b019022ffd208932f036022ffd208c70b018),
    .INIT_66(256'h022ffd2086b2f03d022ffd11c010b01b022ffd14c002f03c022ffd0d5040b01a),
    .INIT_67(256'h022ffd208d52f03f022ffd208d70b01d022ffd250002f03e022ffd208910b01c),
    .INIT_68(256'h022ffd09c0c1d001022ffd2b03c323a9022ffd2b80c1d000022ffd208930b001),
    .INIT_69(256'h022ffd2086b1d003022ffd09c0c323b1022ffd2b02c1d002022ffd2086b323ad),
    .INIT_6A(256'h022ffd2b00c20be5022ffd2086b20a7a022ffd09c0c20b91022ffd2b01c323b5),
    .INIT_6B(256'h022ffd2500020be5022ffd2089120a81022ffd2086b20b94022ffd09c0c223b8),
    .INIT_6C(256'h022ffd208df20be5022ffd208df20a8b022ffd208df20b97022ffd208df223b8),
    .INIT_6D(256'h022ffd208df20be5022ffd208df20a97022ffd208df20b9a022ffd208df223b8),
    .INIT_6E(256'h022ffd369c00b017022ffd1d0001c010022ffd0b0320b134022ffd250000b016),
    .INIT_6F(256'h022ffd208910b136022ffd208d30b018022ffd208cd1e010022ffd208b50b135),
    .INIT_70(256'h022ffd208b11e010022ffd208c70b13b022ffd208b50b019022ffd250001e010),
    .INIT_71(256'h022ffd1d0000b01b022ffd0b0321e010022ffd250000b13c022ffd208910b01a),
    .INIT_72(256'h022ffd208b70b13e022ffd208cb0b01c022ffd208b91e010022ffd369cd0b13d),
    .INIT_73(256'h022ffd208b51e010022ffd208b90b13f022ffd250000b01d022ffd208911e010),
    .INIT_74(256'h022ffd208cf323dd022ffd2099e1d800022ffd2089119801022ffd208b5363f1),
    .INIT_75(256'h022ffd141061d001022ffd0b113323a9022ffd208931d000022ffd208b10b001),
    .INIT_76(256'h022ffd0b00f1d003022ffd14106323b1022ffd141061d002022ffd14106323ad),
    .INIT_77(256'h022ffd2086a20d85022ffd0b00e2f013022ffd2086a0b001022ffd04010323b5),
    .INIT_78(256'h022ffd2086a2f013022ffd0b00c0b001022ffd2086a2f01f022ffd0b00d01004),
    .INIT_79(256'h022ffd2089320891022ffd208b1323e8022ffd208c71d002022ffd208910b032),
    .INIT_7A(256'h022ffd1410632711022ffd0b1131d001022ffd2086a0b032022ffd0100020941),
    .INIT_7B(256'h022ffd2086a20902022ffd0401001004022ffd0b01232711022ffd141061d002),
    .INIT_7C(256'h022ffd2086a2f03a022ffd0b01011001022ffd2086a0b03a022ffd0b01122008),
    .INIT_7D(256'h022ffd1dcff1f000022ffd0bc170b017022ffd250001d000022ffd208910b016),
    .INIT_7E(256'h022ffd34a3a1f000022ffd1dcff0b019022ffd0bc161f000022ffd34a340b018),
    .INIT_7F(256'h022ffd0bc181f00002bff334a340b01b02bff01dcff1f000022ffd0bc190b01a),
    .INITP_00(256'h35e369d73199ba33836b7fc3333f8dad690b2b5a948a2eb853819d896c19bf39),
    .INITP_01(256'ha7c4148c999c742305871345b50c12fa85120c638923baa14a23aa8d25a59917),
    .INITP_02(256'hde7764d2950bb1379764dbe89a990509d93b9eea35b681ab44049f185616b9b8),
    .INITP_03(256'h6a15a803c152cfd6eb4690b68d40f35f0919ecd60423cd5e148e427b190fde1d),
    .INITP_04(256'hac21e8b9043cf9af9d1eb5413396254974355de261a77116aa27371dba86f067),
    .INITP_05(256'h050aaced647532b82bae23789b1f9409b13e03b99dbff278e505b907e872c77b),
    .INITP_06(256'h211f060c3f02998a56aab2a5132ac697131a7f5e2bef6ff52f47b9aaa4bf3850),
    .INITP_07(256'h63da8e77e66d917b9ca33e33a1e5e9dd8bbb2e0132372ecd0a133c9d1fbdf564),
    .INITP_08(256'h7c17292b04080380701e899c1e0198ebe59a9297bd9d4a28013fa830e5139a1b),
    .INITP_09(256'h09a4fb490088a132204e2fa8989f046a1f03874ee5fbf616da99a8b1a814795a),
    .INITP_0A(256'h178690e2f8d6c08eb11dc04e4c6b6c5736ede0f99237b085bd312975992e2c2b),
    .INITP_0B(256'h98b82fb50a86aa37bf7d22b0ba6867cc4cdba6a4126b605b5f859019de6ec0e1),
    .INITP_0C(256'h5bcceb69e7d04df8e8edf95767686346ec52f2d6f7d84ce4556350c445012a05),
    .INITP_0D(256'h6cd5466944c8fa6543c3cc4143cbce4176f2f7d95cf355d4724bcee450c37279),
    .INITP_0E(256'h66fe7c75ff627f6a79d36bfd4d4276f4fb6a64f8f3507adacaeb606ae7d66f76),
    .INITP_0F(256'heac2687964cef07241617eeb7d657efbe57aed7feb4679fdee71cde7736af273),
