    .INIT_00(256'h032c2b20b9a2002001d0d1226052ff00032c1620a8b01f0001d0d020b9728000),
    .INIT_01(256'h020c492b6c9209020001e02b00a01001020c49208912004c0001f020a9720033),
    .INIT_02(256'h020c4909d081d0020001c009e0832060020c4909f081d0010001d00125d208f3),
    .INIT_03(256'h02f12c2086b1d01002f12a00cd03249402f1282086b1d00000110009c0832256),
    .INIT_04(256'h02f12d2086b1d00802f12b00cf03271102f1292086b1d00402f12e00ce03265f),
    .INIT_05(256'h020c4920b08010600001f03660932426025000192011d08202f12f20891327bb),
    .INIT_06(256'h020c4922008208bf0001d02093020902020c49208910109f0001e02261a208f6),
    .INIT_07(256'h02f62a2023b22ffd02f7282023220891020c4920891208d70001c0208cd208c7),
    .INIT_08(256'h001500202440b000001400326283202f02f42e1d0020d08002f52c0b00209002),
    .INIT_09(256'h02f62b2024d011ff02f72932628010ff0017001d0033602f0016000b0020d001),
    .INIT_0A(256'h0001f0209301b200022c15209021b10002f42f010021900102f52d20b080121f),
    .INIT_0B(256'h0001d02023b09001020c49202322f0000001e02089101001020c49220083e029),
    .INIT_0C(256'h000170202442b000020c4932638250000001c01d0023202f020c490b0020d040),
    .INIT_0D(256'h0001602024d010ff0037f0326382bfff02f1291d0032bf7e00310f0b0022b00c),
    .INIT_0E(256'h000150010010300f0036f02f01e0900102f12b010002d01100310f20b082d010),
    .INIT_0F(256'h00014020897360420035f0208b70d02002f12d2091e0900d00310f2f0322d001),
    .INIT_10(256'h00110020893090060034f0208cb0900602f12f226c52203d00310f2089309006),
    .INIT_11(256'h02f12e2087c0900702f12c208723604902f12a208720d08002f1280bc330900d),
    .INIT_12(256'h0141000bc0a250000144002086b090070141000bc0b09007022c15208e522044),
    .INIT_13(256'h0141000bc08208950146002086b208c90141000bc09208b90145002086b208d5),
    .INIT_14(256'h01410020891208d30144002086b208d70141000bc07208c70147002086b208d9),
    .INIT_15(256'h01410020b342089b0146003265b208db0141000d0082089501450009002208b1),
    .INIT_16(256'h00b8280100025000000170220082089102500020902208990147000101020895),
    .INIT_17(256'h020d250ba0725000020d07220083e05d020cfb209301900100b9292090201019),
    .INIT_18(256'h014b000be0b0900d014a0e0bd0a201ab00ba250bc09201c5001b000bb08201bd),
    .INIT_19(256'h014a001d00c20a53014b000300f20a4c014a00000f03206300ba260bf330d001),
    .INIT_1A(256'h00b217226c020b8b014b003266c20b60014a000d00801101014b003266c01080),
    .INIT_1B(256'h014b002085001000014a002f0140110002f2170301f360660062b0000a01dc93),
    .INIT_1C(256'h014b000307f0311e014a00000b0001e0014b002085020e5f014a002085020b77),
    .INIT_1D(256'h014b000b033000d0014a002f01522017014b003e6c032077014a001d05d1d112),
    .INIT_1E(256'h014a000d008030f8014b003267d14008014a001d00c1410a00ba270300f001e0),
    .INIT_1F(256'h00b2160300332085014b001400e1d048014a00000e032085014b00326861d058),
    .INIT_20(256'h00b82a366c0320880001601c0101d00002fb160b11332088006b202f0131d088),
    .INIT_21(256'h020d25030032208d020d070b0332f002020cfb366950100200b92b2085022017),
    .INIT_22(256'h014b00366c001004014a0e1c0102208d00ba250b1132f002001b002f01301003),
    .INIT_23(256'h014a002fe0e2f239014b002fd0d01220014a002fc0c201a700ba26208502f002),
    .INIT_24(256'h00b219326c02f03a014b001df0101000014a0003f072f201014b002ff0f01203),
    .INIT_25(256'h014b002fd11201d0014a002fc10201b702f21903e032f0240062b0226a401001),
    .INIT_26(256'h014b000b20601100014a000b10520b8b014b000b004201f8014a002fe12201d9),
    .INIT_27(256'h014b003e6c001010014a001ae20201f8014b001ad1020b77014a0018c0001010),
    .INIT_28(256'h014a002f40f01010014b000340701100014a000b40f201e200ba2720e7a01100),
    .INIT_29(256'h00b2181d00120a5c014b00326ad20a56014a001d00020a59014b000b01320b77),
    .INIT_2A(256'h00b82c1d00320bd5000150326b72b02e02fb181d00220bd5006b20326b22b02e),
    .INIT_2B(256'h020d252083520a4c020d0720a7a20b02020cfb20b9120a4c00b92d326bc20b34),
    .INIT_2C(256'h014b0020a8120b8b014a0e20b9420b6000ba25226c001101001b0020ba601080),
    .INIT_2D(256'h014a0020b9720b42014b00226c020b77014a0020bb00100400ba262083501100),
    .INIT_2E(256'h00b21b226c020a4c014b0020bbb201d9014a002083520b42014b0020a8b201d0),
    .INIT_2F(256'h014b0020bc620b8b014a0020835201f802f21b20a9720a4c0062b020b9a20b02),
    .INIT_30(256'h014b0020930010c0014a002090220b77014b000100001014014a0020b0801100),
    .INIT_31(256'h014b003625c01014014a000d00820b42014b000901120b60014a002200801101),
    .INIT_32(256'h014a000d04001014014b00362c901100014a000d080201e200ba270900e01100),
    .INIT_33(256'h00b21a0d01020b42014b00362c320a59014a000d02020b42014b00362c620b77),
    .INIT_34(256'h00b82e326db010020001400d00420a5c02fb1a0900e20b42006b20362c020a56),
    .INIT_35(256'h020d250300f2d00f020d072b04e01002020cfb2f03320bd900b92f090162d00f),
    .INIT_36(256'h014b000900d32145014a0e226c51d00200ba25326ef0b002001b001d00e20bd9),
    .INIT_37(256'h014a001d04920a4c014b000900620b02014a00366c520a4c00ba260d02020b34),
    .INIT_38(256'h00b21d208d501101014b00366c501080014a001d05320a4c014b00326ef20b02),
    .INIT_39(256'h014b002093901008014a00013000110002f21d0b20220b8b0062b02089120b60),
    .INIT_3A(256'h014b00208b720b48014a00366e7201d0014b001c32020b48014a001130120b77),
    .INIT_3B(256'h014b00208c120a4c014a00226c520b02014b002089320a4c014a0020897201d9),
    .INIT_3C(256'h014a000b00220b8b014b002020c201f8014a002020320a4c00ba272089120b02),
    .INIT_3D(256'h00b21c0b002010c0014b002021520b77014a00326fb01018014b001d00201100),
    .INIT_3E(256'h001a0020b08010180250002021e20b4802fb1c326fb20b60006b201d00301101),
    .INIT_3F(256'h00d8ff0b00201018014a002020c0110000d1ff20203201e2001b002270a01100),
    .INIT_40(256'h00daff0b00220b48014a002021520a5900d9ff3270720b48014a001d00220b77),
    .INIT_41(256'h00020020b08010020250002021e20a5c02fb253270720b48014b001d00320a56),
    .INIT_42(256'h014a042f0322d010014a00010000100200d1ff208f620bdd001a00010602d010),
    .INIT_43(256'h014a042093032145014a04209021d003014a04010000b002014a042d00320bdd),
    .INIT_44(256'h0022a03677620a4c014a041d00120b02014a040b01e20a4c014a042200820b34),
    .INIT_45(256'h02500020d4920a4c02f2260b51720b020062b00b41620a4c020d180120020b02),
    .INIT_46(256'h014b000b41820b8b014a060421020b60000b902f91701101000a802f81601080),
    .INIT_47(256'h014b002f91920b52014a062f81820b77014b0020d490100c014a060b51901100),
    .INIT_48(256'h014b0020d4920a4c014a060b51b201d9014b000b41a20b52014a0604210201d0),
    .INIT_49(256'h001a000b41c20a4c0003800421020b020002102f91b20a4c0250002f81a20b02),
    .INIT_4A(256'h00d2ff2f91d20b8b0033012f81c201f80032aa20d4920a4c001b000b51d20b02),
    .INIT_4B(256'h00daff01202010c0014a003273a20b7700d3ff0d2020101c014a000421001100),
    .INIT_4C(256'h001a00209c60101c000380209b920b52000210209ce20b60014b082f21e01101),
    .INIT_4D(256'h014a00208f00101c00d2ff326fd011000033021d001201e20032cc0b03201100),
    .INIT_4E(256'h014b082f21e20b5200daff0120420a59014a00227b720b5200d3ff0502020b77),
    .INIT_4F(256'h0032f02f01401002001a000b11720a5c0003800b01620b5200021020f5620a56),
    .INIT_50(256'h00d3ff348352d011014a001f1ff0100200d2ff1d0ff20be10033042f1152d011),
    .INIT_51(256'h02fb272f115201b1014b082f014201a700daff0b11920b34014a000b01820be1),
    .INIT_52(256'h00100c0b01a0110000084034835010100009501f1ff201f80250001d0ff20a4c),
    .INIT_53(256'h0131001d0ff20b770148082f1150101001490e2f014011000011000b11b201ed),
    .INIT_54(256'h036d570b11d0110001d1000b01c01014036d4d34835201f80190011f1ff20b42),
    .INIT_55(256'h00d5081f1ff20b770250001d0ff010140018ff2f115011000019ff2f014201ed),
    .INIT_56(256'h0018ff3676c20b480019ff1d0003216e0011020b0321d002036d5d348350b002),
    .INIT_57(256'h0001501d001201ed03ed6a327650110001d1031d000010180250000b013201f8),
    .INIT_58(256'h01410e1d0030b0020118013276920b770018ff1d002010180000403276701100),
    .INIT_59(256'h00190b20bb0201f80118082276c20b5203ed6220ba63216e0140083276b1d003),
    .INIT_5A(256'h00084020bc6011000009502276c201ed02500020bbb011000011042276c0101c),
    .INIT_5B(256'h001102209c62b04e03ed73209f6201a701b905209b920b77019818209ce0101c),
    .INIT_5C(256'h000180208f032195025000326fd1d0010018ff1d0010300f0019ff0b03209001),
    .INIT_5D(256'h0141063678320b080149001d00832186014106227b70d00200381f030df09002),
    .INIT_5E(256'h001102208912b04f014900208b52b80f014106208d32b40f014900208b52b20f),
    .INIT_5F(256'h03ad82326fd2d01001d8141d001010e0036d800b0322b10f01d90b2099e2b08f),
    .INIT_60(256'h03ad801d0102090201d808227b701002025000050202d010001104208f00101c),
    .INIT_61(256'h00b20c208df2020c020e5f208d920203037001208b1220080250003679020930),
    .INIT_62(256'h0005401d0012021500ba0f0b0323219000b40e2099e1d00200b30d208910b002),
    .INIT_63(256'h0006a0227b72021e01450e050203219001450e208f01d003003403326fd0b002),
    .INIT_64(256'h01470e208d92093001470e208b1209020007a03679d010000036071d02020b08),
    .INIT_65(256'h001d000b0322b40f0037032099e2b20f01470e2089120b0801470e208df22008),
    .INIT_66(256'h032dc1030df2b10f01d602208f02b08f000820326fd2b04f001e001d0012b80f),
    .INIT_67(256'h032e1f208b12d01001d604367aa0101c032de91d0402d01001d603227b7010e0),
    .INIT_68(256'h036da62099e208b701cd30208912091e001a00208df2f032001900208d901001),
    .INIT_69(256'h0108f0208f0208cd009f08326fd226c5032dad1d0012089301ce400b03220897),
    .INIT_6A(256'h013e0036017208c1011d011d08025000013a00227b720891013900030df208c5),
    .INIT_6B(256'h00bf31208912089300be30208c9208cf001d00208cd208b1022da2208d3208b5),
    .INIT_6C(256'h0129f0326fd208c10108e01d001208cb032db70b032208c101cd502099e25000),
    .INIT_6D(256'h02f810208f6208d3022db0227b725000011d01030df20893013a00208f0208d7),
    .INIT_6E(256'h0140060b01e2089300b01322008208c5003a0320902208b302f91101008208b7),
    .INIT_6F(256'h037000208f02089302fa12327bf208d5004a00367db208bb0140061d00425000),
    .INIT_70(256'h00b237030bf2089100be31208f02086a00bd30227c40300f0250000504009001),
    .INIT_71(256'h01cf200b01f20893001f002f03b208bb001a000b00e208b1001900208f625000),
    .INIT_72(256'h013a002023b1400e0129e0202321400e0108d0367d703008032dce1900109002),
    .INIT_73(256'h00b23c2024425000001f00327d420891022dc71d0022086a011f010b0021400e),
    .INIT_74(256'h0139002024d01f00010820327d420b60032dd71d0030110001cf500b002010c0),
    .INIT_75(256'h001f002f01f20b8e022dd02280501c00011f010100201d01013a0020b0801e00),
    .INIT_76(256'h0139001d00220b600118022200801100032ddf20918010a001cf300108225000),
    .INIT_77(256'h02f8101d01001c00022dd8327f601d00011f011d00801e00013800327f601f00),
    .INIT_78(256'h014006208f003f8100b013367e820b7e003a031d0202500002f911327f620b8e),
    .INIT_79(256'h0370002280505f0002fa120100203c3f004a00208f603d7c0140060504003e3c),
    .INIT_7A(256'h00b237030bf20b8e00be31208f005c0000bd30367ef05d030250001d04005e40),
    .INIT_7B(256'h001f001d08003e7f001a002280503fff0019000100220b7e001800208f625000),
    .INIT_7C(256'h0129e0208f605e800108d0030bf05f00032df7208f003cff01cf203601703dfd),
    .INIT_7D(256'h00bf392020c25000022df02020320b8e011f012280505c00013a000100205d00),
    .INIT_7E(256'h001f002021525000032e043280020b6001df001d00201101003ff00b002010c0),
    .INIT_7F(256'h0108202021e03dfe032e043280003eff01df021d00303fff00b23c0b00220b7e),
    .INITP_00(256'h78e7cea77da1561c69275366c07e70fc61c4d902da9078a4e81e5b2ef2916c99),
    .INITP_01(256'ha1a042118a22c231951ac71033493fcc966f3d6e97ee7a517367089414317040),
    .INITP_02(256'h74d15130339cf20ba7878a10971b0f1008ae19a9049488ca597dead73f2b5f1f),
    .INITP_03(256'h26a6073c3ba783ae1c3583af192380b8903d752d122225b802ba97bf2c2da880),
    .INITP_04(256'h82882d99ae8817922728613d94340c0983babea9a78f1a255b6c41152885c2b1),
    .INITP_05(256'hb694eebf1b9506b3a7bcba9ca99a0b27d053c2a0b4aceb9b1e3601801e1f1293),
    .INITP_06(256'habbd00b5b033b214d3fe440bbc31dd280119309c988e14a9b6b2ba058a3f0d8f),
    .INITP_07(256'h38960c31b5c2f4929aaa2c3c36278b0da68002bb8a920e1c8dbf702093ab3305),
    .INITP_08(256'h09090e24bc168a356f6813f787a412a80880873106b011ad3fc0c330151eb419),
    .INITP_09(256'h8eb7871207b39a3312303f1f8e363f192f872e8cb0a71728242aaed99f30ad06),
    .INITP_0A(256'hb15c3ce40bbb03ff0fd79d99ff1744180f8a811d1a1b94c867bb3dadae111eac),
    .INITP_0B(256'h7435cba01f3529aab18d3a8296f68a951d68952b9907eabeac17699c99281184),
    .INITP_0C(256'he8b27f9ec136b6003b2ba9939f3aa5ba8fb434073b023ca70def5b5761805b2f),
    .INITP_0D(256'h49671281a708a7674d7108babfa75410348d97e104a3a2a38a0b488ecea53fb7),
    .INITP_0E(256'h51c2b785a508643804d1992888b9f91da1bb759f29ad97783a028c2804a735ec),
    .INITP_0F(256'h2f532ab2b64503a4b7491b932c82c8958482831f09baa1747be3ab3f18b91b51),
