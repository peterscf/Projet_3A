    .INIT_00(256'h0000000b2181daa000000014b003241000000014a001fb0200000014b001da80),
    .INIT_01(256'h0000000b82c1fb02000000001501dac00000002fb183241000000006b201fb02),
    .INIT_02(256'h00000020a813241000000020a631fb0300000020a571da000000000b92d32410),
    .INIT_03(256'h00000014b002242200000014a0e324100000000ba251fb0300000001b001dae0),
    .INIT_04(256'h00000014a00001b000000014b00000a000000014a00208c60000000ba262070b),
    .INIT_05(256'h0000000b21b00bc000000014b002091400000014a00208e700000014b0020904),
    .INIT_06(256'h00000014b00206e500000014a0000ce00000002f21b206e5000000062b000cf0),
    .INIT_07(256'h00000014b00206e500000014a0000cb000000014b00206e500000014a0000cd0),
    .INIT_08(256'h00000014b00207aa00000014a002070b00000014b002242200000014a00208d5),
    .INIT_09(256'h00000014a00208c600000014b002070b00000014a00207470000000ba2722008),
    .INIT_0A(256'h0000000b21a2b40f00000014b002b20f00000014a00208d500000014b002011d),
    .INIT_0B(256'h0000000b82e207aa000000001402077c0000002fb1a0100200000006b202b80f),
    .INIT_0C(256'h00000020a812011d00000020a63208c600000020a572070b0000000b92f22008),
    .INIT_0D(256'h00000014b002b80f00000014a0e2b40f0000000ba252b20f00000001b00208d5),
    .INIT_0E(256'h00000014a002f03200000014b000100100000014a002f01e0000000ba2601000),
    .INIT_0F(256'h0000000b21d2070d00000014b002071100000014a002073100000014b0020798),
    .INIT_10(256'h00000014b002b20f00000014a00208c60000002f21d2070b000000062b0224b4),
    .INIT_11(256'h00000014b002f03200000014a000100200000014b002b80f00000014a002b40f),
    .INIT_12(256'h00000014b002070d00000014a002074500000014b00224f500000014a0020798),
    .INIT_13(256'h00000014a00206f600000014b00206ec00000014a00206ec0000000ba270bc33),
    .INIT_14(256'h0000000b21c0bc0a00000014b00206e500000014a000bc0b00000014b002075f),
    .INIT_15(256'h00000001a000bc0800000025000206e50000002fb1c0bc0900000006b20206e5),
    .INIT_16(256'h0000000d8ff2070b00000014a00206e50000000d1ff0bc0700000001b00206e5),
    .INIT_17(256'h0000000daff208c600000014a00324630000000d9ff0d00800000014a0009002),
    .INIT_18(256'h000000002000100000000025000220080000002fb252077c00000014b0001010),
    .INIT_19(256'h00000014a040ba0700000014a00220080000000d1ff207aa00000001a002077c),
    .INIT_1A(256'h00000014a040be0b00000014a040bd0a00000014a040bc0900000014a040bb08),
    .INIT_1B(256'h000000022a01d00c00000014a040300f00000014a04000f000000014a040bf33),
    .INIT_1C(256'h00000025000224af0000002f22632474000000062b00d00800000020a7432474),
    .INIT_1D(256'h00000014b00206ca00000014a062f01400000000b900301f00000000a80000a0),
    .INIT_1E(256'h00000014b000307f00000014a06000b000000014b00206ca00000014a06206ca),
    .INIT_1F(256'h00000014b000b03300000014a062f01500000014b003e4af00000014a061d05d),
    .INIT_20(256'h00000001a000d0080000000038032485000000002101d00c000000250000300f),
    .INIT_21(256'h0000000d2ff03003000000033011400e000000032aa000e000000001b003248e),
    .INIT_22(256'h0000000daff364af00000014a001c0100000000d3ff0b10200000014a002f013),
    .INIT_23(256'h00000001a0003003000000003800b033000000002103649d00000014b08206ca),
    .INIT_24(256'h00000014a00364af0000000d2ff1c010000000033020b102000000032cc2f013),
    .INIT_25(256'h00000014b082fe0e0000000daff2fd0d00000014a002fc0c0000000d3ff206ca),
    .INIT_26(256'h000000032f0324af00000001a001df010000000038003f07000000002102ff0f),
    .INIT_27(256'h0000000d3ff2fd1100000014a002fc100000000d2ff03e0300000003304224ac),
    .INIT_28(256'h0000002fb270b20600000014b080b1050000000daff0b00400000014a002fe12),
    .INIT_29(256'h0000000100c3e4af000000008401ae20000000009501ad100000002500018c00),
    .INIT_2A(256'h000000131002f40f00000014808034070000001490e0b40f0000000110020bd6),
    .INIT_2B(256'h00000036ab3208d50000001d1002092e00000036aa9206af000000190012092a),
    .INIT_2C(256'h0000000d5082200800000025000207aa000000018ff2077c000000019ff01000),
    .INIT_2D(256'h000000018ff0d020000000019ff36171000000011020d04000000036ab90900f),
    .INIT_2E(256'h000000001500900e0000003eac63616c0000001d1030d0800000002500036171),
    .INIT_2F(256'h0000001410e36165000000118010d040000000018ff36168000000000400d080),
    .INIT_30(256'h0000000190b3615f000000118080d0100000003eabe36162000000140080d020),
    .INIT_31(256'h000000008400901600000000950324ce000000250000d004000000011040900e),
    .INIT_32(256'h000000011021d00e0000003eacf0300f0000001b9052b04e000000198182f033),
    .INIT_33(256'h000000001800d020000000250000900d000000018ff224b4000000019ff324dd),
    .INIT_34(256'h00000014106324dd000000149001d04900000014106090060000000381f364b4),
    .INIT_35(256'h000000011022070b000000149002074f00000014106364b4000000149001d053),
    .INIT_36(256'h0000003aade2070d0000001d8142071100000036adc207310000001d90b207b3),
    .INIT_37(256'h0000003aadc208c60000001d8082070b000000250002073b00000001104224b4),
    .INIT_38(256'h0000000b20c2f03200000020bbb0100000000037001208d50000002500020113),
    .INIT_39(256'h00000000540207aa0000000ba0f2077c0000000b40e010000000000b30d2d003),
    .INIT_3A(256'h000000006a0208d50000001450e201130000001450e208c60000000340322008),
    .INIT_3B(256'h0000001470e2f0320000001470e01000000000007a0207700000000360701060),
    .INIT_3C(256'h00000001d00207aa000000037032077c0000001470e010000000001470e2d003),
    .INIT_3D(256'h00000032b1d01f000000001d60201e000000000082001d0000000001e0022008),
    .INIT_3E(256'h00000032b7b01d010000001d6042ff1200000032b452fe110000001d6032fd10),
    .INIT_3F(256'h00000036b021d0ff0000001cd300b00f00000001a0020bd6000000019002fd1e),
    .INIT_40(256'h000000108f02f00f00000009f080300700000032b090b00f0000001ce4032507),
    .INIT_41(256'h00000013e000900e00000011d012219300000013a0020941000000139002092a),
    .INIT_42(256'h0000000bf312f00b0000000be300901b00000001d003251000000022afe0d004),
    .INIT_43(256'h000000129f032522000000108e01d00e00000032b130300f0000001cd502b04e),
    .INIT_44(256'h0000002f8100bd1000000022b0c0b20600000011d010b10500000013a000b004),
    .INIT_45(256'h000000140061cd000000000b00203f0100000003a030bf120000002f9110be11),
    .INIT_46(256'h0000003700011d010000002fa123252200000004a001ef20000000140061ee10),
    .INIT_47(256'h0000000b2372fe110000000be312fd100000000bd3013f000000002500013e00),
    .INIT_48(256'h0000001cf202011300000001f00208c600000001a00224fb000000019002ff12),
    .INIT_49(256'h00000013a0001000000000129e02d103000000108d00100000000032b2a208d5),
    .INIT_4A(256'h0000000b23c0b01e00000001f002200800000022b23207aa00000011f012077c),
    .INIT_4B(256'h000000139000b416000000108200120000000032b33365850000001cf501d001),
    .INIT_4C(256'h00000001f002f91700000022b2c2f81600000011f0120aa500000013a000b517),
    .INIT_4D(256'h0000001390020aa5000000118020b51900000032b3b0b4180000001cf3004210),
    .INIT_4E(256'h0000002f8100b41a00000022b340421000000011f012f919000000138002f818),
    .INIT_4F(256'h000000140062f91b0000000b0022f81a00000003a0320aa50000002f9110b51b),
    .INIT_50(256'h0000003700020aa50000002fa120b51d00000004a000b41c0000001400604210),
    .INIT_51(256'h0000000b2370d2020000000be31042100000000bd302f91d000000250002f81c),
    .INIT_52(256'h00000001f002084800000001a002f21e00000001900012020000000180032556),
    .INIT_53(256'h000000129e01d001000000108d00b03200000032b53208400000001cf2020833),
    .INIT_54(256'h0000000bf392076a00000022b4c3250700000011f011d00200000013a00324e9),
    .INIT_55(256'h00000001f002f21e00000032b60012040000001df00225c600000003ff005020),
    .INIT_56(256'h000000108202f01400000032b600b1170000001df020b0160000000b23c20cb2),
    .INIT_57(256'h00000022b59346af00000011f011f1ff00000013a001d0ff000000139002f115),
    .INIT_58(256'h00000032b692f1150000001cf502f0140000000b2380b11900000001f000b018),
    .INIT_59(256'h00000011f010b01a00000013a00346af000000139001f1ff000000108201d0ff),
    .INIT_5A(256'h00000032b711d0ff0000001cf302f11500000001f002f01400000022b620b11b),
    .INIT_5B(256'h00000011f010b11d000000138000b01c00000013900346af000000118011f1ff),
    .INIT_5C(256'h00000003a031f1ff0000002f9111d0ff0000002f8102f11500000022b6a2f014),
    .INIT_5D(256'h00000004a0036579000000140061d000000000140060b0320000000b002346af),
    .INIT_5E(256'h0000000bd3020870000000250002083300000037000208480000002fa122092e),
    .INIT_5F(256'h00000001900324e9000000018001d0010000000b2370b0320000000be3120840),
    .INIT_60(256'h00000032b89030df0000001cf202076a00000001f003250700000001a001d002),
    .INIT_61(256'h00000011f012072f00000013a0036592000000129e01d008000000108d0225c6),
    .INIT_62(256'h0000001df002081800000003ff02070b0000000bf392072f00000022b822074d),
    .INIT_63(256'h0000001df022076a0000000b23c324e900000001f001d00100000032b960b032),
    .INIT_64(256'h00000013a003659f000000139001d01000000010820225c600000032b9605020),
    .INIT_65(256'h0000000b2382070b00000001f002075900000022b8f2075300000011f012072b),
    .INIT_66(256'h00000010820324e900000032ba01d0010000001cf000b0320000000b03720818),
    .INIT_67(256'h00000022b981d02000000011f01225c600000013a0005020000000139002076a),
    .INIT_68(256'h00000032ba9207590000001cf50207530000000b2032072b00000001f00365ac),
    .INIT_69(256'h00000011f011d00100000013a000b0320000001390020818000000108202070b),
    .INIT_6A(256'h00000032bb1225c60000001cf30030df00000001f002076a00000022ba2324e9),
    .INIT_6B(256'h00000011f0120753000000138002072b00000013900365b9000000118011d040),
    .INIT_6C(256'h00000003a030b0320000002f911208180000002f8102070b00000022baa20759),
    .INIT_6D(256'h00000004a00030df000000140062076a00000014006324e90000000b0021d001),
    .INIT_6E(256'h00000020bcf2074d0000002500036017000000370001d0800000002fa12225c6),
    .INIT_6F(256'h0000000960820818000000095082070b0000002f503207430000000950820747),
    .INIT_70(256'h000000096082076a00000009508324e90000002f6051d0010000002f5040b032),
    .INIT_71(256'h000000096080100800000009508207700000002f631225c60000002f530030df),
    .INIT_72(256'h000000096081d004000000095080b01e0000002f638220080000002f5372077c),
    .INIT_73(256'h000000015ef3261f000000250000d0040000002f606090020000002f53c36634),
    .INIT_74(256'h0000002d60a01e400000002d50901f0a000000011002069e0000000160720678),
    .INIT_75(256'h00000020bbb09d070000003700120658000000250000120b0000002d10b011b3),
    .INIT_76(256'h0000002f8341ce100000000ba122dd080000000b9112de090000000b8102df0a),
    .INIT_77(256'h0000000bd37225e300000001200365e00000002fa361cf200000002f935365e0),
    .INIT_78(256'h0000001a9400b01600000018830225d60000000b43113f000000000b33011e01),
    .INIT_79(256'h0000002f8341d0ff000000112012f1150000003abed2f0140000001ba000b117),
    .INIT_7A(256'h00000032c19012000000001c2d0206600000002fa36325ef0000002f9351f1ff),
    .INIT_7B(256'h0000000ba360b0180000000b9352f2200000000b8341420000000022be20d0ff),
    .INIT_7C(256'h000000094081d0ff000000013002f115000000012002f0140000002f20f0b119),
    .INIT_7D(256'h0000001b90001200000000188402066000000032cab325fb0000001d4011f1ff),
    .INIT_7E(256'h000000133000b01a000000112012f2210000003ac00142000000001ba000d0ff),
    .INIT_7F(256'h00000022bf31d0ff0000002fa362f1150000002f9352f0140000002f8340b11b),
    .INITP_00(256'h3d913d103d13189c16278bae82258225278e3c91821396309c01163e1eb70135),
    .INITP_01(256'h9d329b3a11321aad3611340b071316bc99100e2a12a90d32823990a6bc1a270d),
    .INITP_02(256'h269a37021a1e0f18a8bc9021963d8b3d91b99aaa3a15a9193217360ba9829b04),
    .INITP_03(256'hb29c3e022d083094301f1226288f1201351a98909919121d97839ab736210a38),
    .INITP_04(256'h2f001518b5be39373d2208b2089c0f31a2b4b4adac1ebd1805141d9331b1bea4),
    .INITP_05(256'h34288e3e9f2132229aa00720bc3d91b22ba9293f18b7018c3b0db0bf9a22b68b),
    .INITP_06(256'h19aebb9a19ba03840510a606370da237182701311eab81918aa4371bb02d9886),
    .INITP_07(256'h3a1a2dabb014a4020497b88318bea8b82ba80c00318b1c28383588bb1120b6b7),
    .INITP_08(256'h10140e25b5b8b81881a1892f963daa349b9097bbac0c1e0b80bca5a21f951a3e),
    .INITP_09(256'h86b3073f88ab940aaaaa86be21379939300e839598a02400b495829a26a1ab24),
    .INITP_0A(256'h888a20b70aa00e02372a0985bf9512b29c023d302931bb10050a04acaa3ab816),
    .INITP_0B(256'h36078f148aa1ab22a30017ab14a78e05801eb428b2bbbb110d33b994a18b0939),
    .INITP_0C(256'h0b10aab906b53eb1873e1802202d10b90815a5270313b10e84221892a32bb3a5),
    .INITP_0D(256'h190cb1869cad2825a31d91381e2982830d122e3e35a53b9714342988a98c9020),
    .INITP_0E(256'h148aa42b9532b486a6283fa1860493a2a0372424120f3ea80405b8af89822128),
    .INITP_0F(256'h20b23a8abc228a1c1791182833369b10bbb412b2a9063eba9da4bb9c932d1134),
