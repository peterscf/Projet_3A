    .INIT_00(256'h022ffd206581f000022ffd09d070b01a022ffd206581f000022ffd09e070b019),
    .INIT_01(256'h022ffd206e51f000022ffd00cd00b01c022ffd206e51f000022ffd09c070b01b),
    .INIT_02(256'h022ffd206e5208d5022ffd00cf036017022ffd206e51f000022ffd00ce00b01d),
    .INIT_03(256'h022ffd2070d1d002022ffd20741324b4022ffd2072f1d001022ffd2070b0b032),
    .INIT_04(256'h022ffd14c002f01e022ffd0d50401001022ffd01c0022008022ffd2071732507),
    .INIT_05(256'h022ffd2500011d01022ffd2070b0bf12022ffd206e50be11022ffd11c010bd10),
    .INIT_06(256'h022ffd2b80c2fe11022ffd2070d2fd10022ffd2074f13f00022ffd2075113e00),
    .INIT_07(256'h022ffd2b02c0b00f022ffd206e520bd6022ffd09c0c2ff12022ffd2b03c03f01),
    .INIT_08(256'h022ffd09c0c0307e022ffd2b01c0b03b022ffd206e52f00f022ffd09c0c03007),
    .INIT_09(256'h022ffd206e536243022ffd09c0c1c0e0022ffd2b00c03e7e022ffd206e50be0e),
    .INIT_0A(256'h022ffd207591d000022ffd207590b016022ffd2500020941022ffd2070b2092a),
    .INIT_0B(256'h022ffd207591f000022ffd207590b018022ffd207591f000022ffd207590b017),
    .INIT_0C(256'h022ffd0b0321f000022ffd250000b01a022ffd207591f000022ffd207590b019),
    .INIT_0D(256'h022ffd207471f000022ffd2072f0b01c022ffd3683a1f000022ffd1d0000b01b),
    .INIT_0E(256'h022ffd2072f22243022ffd250003623c022ffd2070b1f000022ffd2074d0b01d),
    .INIT_0F(256'h022ffd25000207bb022ffd2070b2070b022ffd2072b207aa022ffd207412078b),
    .INIT_10(256'h022ffd20733208d5022ffd3684722008022ffd1d0002077c022ffd0b03201004),
    .INIT_11(256'h022ffd2500001002022ffd2070b2b80f022ffd207312b40f022ffd207452b20f),
    .INIT_12(256'h022ffd2070b01000022ffd2072f22008022ffd2072f207aa022ffd207332077c),
    .INIT_13(256'h022ffd2070d3227e022ffd2072b0d004022ffd207490900e022ffd208182f032),
    .INIT_14(256'h022ffd141062f008022ffd1410609018022ffd141062f007022ffd0b11309017),
    .INIT_15(256'h022ffd206e42f00a022ffd040100901a022ffd0b00f2f009022ffd1410609019),
    .INIT_16(256'h022ffd206e42f033022ffd0b00d09016022ffd206e42f00b022ffd0b00e0901b),
    .INIT_17(256'h022ffd2074136264022ffd2070b1d00a022ffd206e40300f022ffd0b00c2b04e),
    .INIT_18(256'h022ffd206e422425022ffd0100032424022ffd2070d0d002022ffd2072b09002),
    .INIT_19(256'h022ffd0b0121d00b022ffd1410622424022ffd1410636267022ffd0b1131d00e),
    .INIT_1A(256'h022ffd206e42dc01022ffd0b01103c0f022ffd206e40bc07022ffd0401036271),
    .INIT_1B(256'h022ffd250002070b022ffd2070b206e5022ffd206e42070d022ffd0b0102074d),
    .INIT_1C(256'h022ffd0bc1620753022ffd348ae36275022ffd1dcff1d00d022ffd0bc1722003),
    .INIT_1D(256'h022ffd1dcff20731022ffd0bc1936279022ffd348b41d00f022ffd1dcff22441),
    .INIT_1E(256'h022ffd348b40d008022ffd1dcff3244a022ffd0bc181d00c022ffd348ae22431),
    .INIT_1F(256'h022ffd0bc1a0d020022ffd348ae0900d022ffd1dcff22422022ffd0bc1b3244a),
    .INIT_20(256'h022ffd1dcff36288022ffd0bc1d1d04f022ffd348b409006022ffd1dcff36424),
    .INIT_21(256'h022ffd348b422425022ffd1dcff32424022ffd0bc1c0d002022ffd348ae09002),
    .INIT_22(256'h022ffd328922070b022ffd1dd002074f022ffd0bd203628f022ffd250001d053),
    .INIT_23(256'h022ffd208ba1d052022ffd0bc1622423022ffd208ae207c2022ffd0bc17207b3),
    .INIT_24(256'h022ffd1dd0009006022ffd0bd2120762022ffd208c02074d022ffd0bc20362a6),
    .INIT_25(256'h022ffd0bc1820762022ffd208ae2070d022ffd0bc1936422022ffd3289b1d020),
    .INIT_26(256'h022ffd0bd2220717022ffd208c036422022ffd0bc211d030022ffd208ba09006),
    .INIT_27(256'h022ffd208ae3a422022ffd0bc1b206d8022ffd328a409006022ffd1dd0020762),
    .INIT_28(256'h022ffd208c02075f022ffd0bc22206f6022ffd208ba00100022ffd0bc1a2d001),
    .INIT_29(256'h022ffd0bc1d362aa022ffd328ad1d055022ffd1dd0022003022ffd0bd232070b),
    .INIT_2A(256'h022ffd0bc23362ae022ffd208ba1d044022ffd0bc1c22441022ffd208ae20753),
    .INIT_2B(256'h022ffd20731362d5022ffd207571d04e022ffd2500022431022ffd208c020731),
    .INIT_2C(256'h022ffd250001d020022ffd2070d09006022ffd206e520762022ffd2070d20745),
    .INIT_2D(256'h022ffd206e5206fb022ffd2070d0120a022ffd207512070d022ffd2072d36422),
    .INIT_2E(256'h022ffd207512fc0a022ffd2072d2fb09022ffd250002fa08022ffd2070b3a422),
    .INIT_2F(256'h022ffd25000206fb022ffd2070d01201022ffd206e52fe33022ffd2070d2fd0b),
    .INIT_30(256'h022ffd206e514a06022ffd2070d14a06022ffd2075514a06022ffd207413a422),
    .INIT_31(256'h022ffd2b00a0bd0a022ffd2b0090bc09022ffd250000bb08022ffd2070b14a06),
    .INIT_32(256'h022ffd01c00206d1022ffd20939206d1022ffd2b08e0bf33022ffd2b1bb0be0b),
    .INIT_33(256'h022ffd01c102fb08022ffd250002fa07022ffd20059206d1022ffd208de206d1),
    .INIT_34(256'h022ffd208de2ff33022ffd01c072fe0b022ffd250002fd0a022ffd208de2fc09),
    .INIT_35(256'h022ffd2500020751022ffd208de36345022ffd01c0d1d054022ffd250002245b),
    .INIT_36(256'h022ffd01c0436422022ffd250001d020022ffd208de09006022ffd01c0120762),
    .INIT_37(256'h022ffd01e003a422022ffd01d00206fb022ffd250000120a022ffd208de2070d),
    .INIT_38(256'h022ffd011002fd0b022ffd010802fc0a022ffd2090d2fb09022ffd01f002fa08),
    .INIT_39(256'h022ffd2b3893a422022ffd25000206fb022ffd208ed01201022ffd209042fe33),
    .INIT_3A(256'h022ffd2093914a06022ffd2b08e14a06022ffd2b63b14a06022ffd2b00a3a422),
    .INIT_3B(256'h022ffd2b37b0bb08022ffd2b00a0ba07022ffd2b1c92fa07022ffd2500014a06),
    .INIT_3C(256'h022ffd2b6490bf33022ffd250000be0b022ffd209390bd0a022ffd2b08e0bc09),
    .INIT_3D(256'h022ffd20939206d1022ffd2b08e206d1022ffd2b5bb206d1022ffd2b62a206d1),
    .INIT_3E(256'h022ffd2bdcb2fd0a022ffd2b10a2fc09022ffd2b6492fb08022ffd250002fa07),
    .INIT_3F(256'h022ffd2b10a2fb3f022ffd2b6c92fa3e022ffd209392ff33022ffd2b08e2fe0b),
    .INIT_40(256'h022ffd2500032305022ffd209390df08022ffd2b08e32325022ffd2bebb1df0c),
    .INIT_41(256'h022ffd2d10836422022ffd2d00818fa0022ffd2b4190ba02022ffd2b00a22422),
    .INIT_42(256'h022ffd2d108206ca022ffd2d008206ca022ffd2b259206ca022ffd2b00a206ca),
    .INIT_43(256'h022ffd2dc082ff0f022ffd2b2892fe0e022ffd2b00a2fd0d022ffd250002fc0c),
    .INIT_44(256'h022ffd250000be11022ffd2df080bd10022ffd2de082070b022ffd2dd0820ae1),
    .INIT_45(256'h022ffd09d0800cf0022ffd09c0820717022ffd2b2892072f022ffd2b00a0bf12),
    .INIT_46(256'h022ffd208e700cd0022ffd25000206e5022ffd09f0800ce0022ffd09e08206e5),
    .INIT_47(256'h022ffd208ed206ec022ffd2090d206ec022ffd250000bc3f022ffd20914206e5),
    .INIT_48(256'h022ffd20904206e5022ffd011000bc3e022ffd010202075f022ffd25000206f6),
    .INIT_49(256'h022ffd0bc0c0ba02022ffd0bd0d206ca022ffd0be0e206ca022ffd0bf0f22422),
    .INIT_4A(256'h022ffd208db206ca022ffd20921206ca022ffd2500036422022ffd2091e18ea0),
    .INIT_4B(256'h022ffd2500003e03022ffd209302fe12022ffd250002fd11022ffd208f32fc10),
    .INIT_4C(256'h022ffd209040be0d022ffd011010bf0c022ffd010802070b022ffd2092120bd6),
    .INIT_4D(256'h022ffd208f900cd0022ffd208d8206e5022ffd208ed0bc0f022ffd208e70bd0e),
    .INIT_4E(256'h022ffd3693900cf0022ffd0d008206e5022ffd0900e00ce0022ffd25000206e5),
    .INIT_4F(256'h022ffd3293d206ec022ffd0d002206ec022ffd0900e0bc3f022ffd25000206e5),
    .INIT_50(256'h022ffd2f116206e5022ffd011000bc3e022ffd370012075f022ffd25000206f6),
    .INIT_51(256'h022ffd2f11a09002022ffd2f11936363022ffd2f1181d058022ffd2f11722422),
    .INIT_52(256'h022ffd010a220762022ffd2f11d20759022ffd2f11c3e363022ffd2f11b0d004),
    .INIT_53(256'h022ffd110012070d022ffd2b00b36422022ffd2b00a1d020022ffd2b6c909006),
    .INIT_54(256'h022ffd1d0ff2070b022ffd209b63a422022ffd2095c206fb022ffd2095701208),
    .INIT_55(256'h022ffd09c082fd3b022ffd250002fc36022ffd370002fb35022ffd3694f2fa34),
    .INIT_56(256'h022ffd250000bf3b022ffd09f080be36022ffd09e080bd35022ffd09d080bc34),
    .INIT_57(256'h022ffd3298720658022ffd1d0d1206a2022ffd3297201b00022ffd1d0d001a01),
    .INIT_58(256'h022ffd209a51d051022ffd001e022422022ffd209a5206e5022ffd001f009c07),
    .INIT_59(256'h022ffd209a509006022ffd001c020762022ffd209a52074b022ffd001d0363c6),
    .INIT_5A(256'h022ffd2f12c0120a022ffd2f12a2070d022ffd2f12836422022ffd011001d020),
    .INIT_5B(256'h022ffd2f12d2fb09022ffd2f12b2fa08022ffd2f1293a422022ffd2f12e206fb),
    .INIT_5C(256'h022ffd209a501201022ffd001f02fe33022ffd250002fd0b022ffd2f12f2fc0a),
    .INIT_5D(256'h022ffd209a514a06022ffd001d014a06022ffd209a53a422022ffd001e0206fb),
    .INIT_5E(256'h022ffd2f62a0bc09022ffd2f7280bb08022ffd209a514a06022ffd001c014a06),
    .INIT_5F(256'h022ffd01500206d1022ffd014000bf33022ffd2f42e0be0b022ffd2f52c0bd0a),
    .INIT_60(256'h022ffd2f62b2fa07022ffd2f729206d1022ffd01700206d1022ffd01600206d1),
    .INIT_61(256'h022ffd001f02fe0b022ffd229712fd0a022ffd2f42f2fc09022ffd2f52d2fb08),
    .INIT_62(256'h022ffd001d00df08022ffd209a53239a022ffd001e01df0c022ffd209a52ff33),
    .INIT_63(256'h022ffd0017018fa0022ffd209a50ba02022ffd001c022422022ffd209a53238e),
    .INIT_64(256'h022ffd00160206ca022ffd037f0206ca022ffd2f129206ca022ffd0310f36422),
    .INIT_65(256'h022ffd001502fe0e022ffd036f02fd0d022ffd2f12b2fc0c022ffd0310f206ca),
    .INIT_66(256'h022ffd00140206ca022ffd035f0206ca022ffd2f12d223b0022ffd0310f2ff0f),
    .INIT_67(256'h022ffd01100206ca022ffd034f036422022ffd2f12f18ea0022ffd0310f0ba02),
    .INIT_68(256'h022ffd2f12e2fe12022ffd2f12c2fd11022ffd2f12a2fc10022ffd2f128206ca),
    .INIT_69(256'h022ffd1410018c00022ffd144000b206022ffd141000b105022ffd229710b004),
    .INIT_6A(256'h022ffd1410020bd6022ffd146003e422022ffd141001ae20022ffd145001ad10),
    .INIT_6B(256'h022ffd14100223b0022ffd144002f40f022ffd1410003407022ffd147000b40f),
    .INIT_6C(256'h022ffd141002b00a022ffd146002070b022ffd141002092a022ffd14500208c6),
    .INIT_6D(256'h022ffd0b82809e08022ffd0017009f08022ffd250000125d022ffd147002b6c9),
    .INIT_6E(256'h022ffd20a8100cd0022ffd20a63206e5022ffd20a5709c08022ffd0b92909d08),
    .INIT_6F(256'h022ffd14b0000cf0022ffd14a0e206e5022ffd0ba2500ce0022ffd01b00206e5),
    .INIT_70(256'h022ffd14a00363b6022ffd14b0019201022ffd14a002070b022ffd0ba26206e5),
    .INIT_71(256'h022ffd0b21736424022ffd14b001d050022ffd14a0022423022ffd14b00208d5),
    .INIT_72(256'h022ffd14b001d020022ffd14a0009006022ffd2f21720762022ffd062b020749),
    .INIT_73(256'h022ffd14b00206fb022ffd14a0001202022ffd14b002070d022ffd14a0036422),
    .INIT_74(256'h022ffd14b00206ca022ffd14a00206ca022ffd14b00206ca022ffd14a003a422),
    .INIT_75(256'h022ffd14a00206ca022ffd14b0036422022ffd14a0018bc0022ffd0ba270bc02),
    .INIT_76(256'h022ffd0b21636410022ffd14b000d040022ffd14a0009002022ffd14b00206ca),
    .INIT_77(256'h022ffd0b82a1da20022ffd0016032410022ffd2fb161fb00022ffd06b201da00),
    .INIT_78(256'h022ffd20a811fb00022ffd20a631da80022ffd20a5732410022ffd0b92b1fb00),
    .INIT_79(256'h022ffd14b0032410022ffd14a0e1fb00022ffd0ba251daa0022ffd01b0032410),
    .INIT_7A(256'h022ffd14a001dae0022ffd14b0032410022ffd14a001fb00022ffd0ba261dac0),
    .INIT_7B(256'h022ffd0b2191fb01022ffd14b001da20022ffd14a0032410022ffd14b001fb00),
    .INIT_7C(256'h022ffd14b0032410022ffd14a001fb01022ffd2f2191da80022ffd062b032410),
    .INIT_7D(256'h022ffd14b001dac0022ffd14a0032410022ffd14b001fb01022ffd14a001daa0),
    .INIT_7E(256'h022ffd14b001fb02022ffd14a001da00022ffd14b0032410022ffd14a001fb01),
    .INIT_7F(256'h022ffd14a003241002bff314b001fb0202bff014a001da20022ffd0ba2732410),
    .INITP_00(256'h5d6650cffac17cf56fcee0c24276fec44cf8ce59635778d978db78d6c076c0f7),
    .INITP_01(256'hee51cb7acff15d727dd468caf0e4f976f9f5f972eaf1f8486b4cccee5b597ed7),
    .INITP_02(256'he3cc7271e66ae2e961e2ef756ff6e84e5cc1f2c1d9cbd7c56c5ec77a5a4644f2),
    .INITP_03(256'hfe7353e97ac3787dcc62ecd479f3507e61556d706d607eedfdf8f6c1f06f5a56),
    .INITP_04(256'h7362f5e94a56fc72e36d607f72c6c2edf4616d6e6d61c0faea4676f4d473ead2),
    .INITP_05(256'he8d3ec497952744cfdd26b55f44871d9cffff04b6b7e63eb76747458ceeafb60),
    .INITP_06(256'hdecd654de7f4d078615fe7f3db667d59e1f3d6cfe66de449d3597a5570d270eb),
    .INITP_07(256'h74da79eee9f875f36df372d3fbfef3666a5dff65e876d2d175e84b6ed8d7eaf5),
    .INITP_08(256'hcef1756c42655e7073d84753f546716ac2d25073fcdfdfc569d462d2efff76d1),
    .INITP_09(256'h737c406546fe5d65c6cd59d16a4fc6fdecfaf5d041e6fd61f054527cf2d07fea),
    .INITP_0A(256'h5fc448c5f0c9efe64cf27bf64e53ddc9d64a595147c252cd404159ddddd07cea),
    .INITP_0B(256'he3d75c646fd855e755794c7554fafecedfd6454c5adaded2cfe65ae64fe25561),
    .INITP_0C(256'h4ef7d07b484156f84653d1e657e55173c2c5fd526e5d7fc4fe64ce79f3584764),
    .INITP_0D(256'h60dd74c1df564bf2c8476778f9c07bdf70e1f6657049f2d765e7e47054cac34b),
    .INITP_0E(256'hd3d0c57c41e2dbe9ca7ccff3e9cae9de69c0e35f755d414bde7d5ef750e6c3f8),
    .INITP_0F(256'h4d4de068fb436edee74dfd456ede524b46ea4d7e4e6e5dfb6e47fb4b4b5e417e),
