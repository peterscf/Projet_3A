    .INIT_00(256'h02f30e012002002000ba36206602ff0000b9353260701f0000b8341f1ff28000),
    .INIT_01(256'h00b50d0b01c2077c00b40c2f2220100102f80c142002004902f20d0d0ff20033),
    .INIT_02(256'h0146082f1151d00200b30e2f0143205d00b70f012001d00100b60e0b11d2076d),
    .INIT_03(256'h014700206601d010014308326143224b0147001f1ff1d0000146081d0ff3212b),
    .INIT_04(256'h0140062f2231d008014006142003252b00b0020d0ff1d00402f70e0120032467),
    .INIT_05(256'h0370000b0200106002f00f2084032212014006208891d0820140062083b325ca),
    .INIT_06(256'h01d40004010207390034f00b1222077c00b439040100109f0250000b12120770),
    .INIT_07(256'h0188402076a22ffd001200326222070b00b43c0401020751032c4f0b12320741),
    .INIT_08(256'h011201030bf0b00003ac2a2076a3202f01ba00226240d08001b9000504009002),
    .INIT_09(256'h01d2020b01f011ff02fa362f03b010ff02f9350b00e3602f02f834207700d001),
    .INIT_0A(256'h00b9352b20f1b20000b834208d51b100022c1f3663019001032c4f190010121f),
    .INIT_0B(256'h019402226550900100b43c010022f00002f20f2b80f0100100ba362b40f3e029),
    .INIT_0C(256'h03ecab220082b00001ba00207922500001b900010823202f0188402f01f0d040),
    .INIT_0D(256'h00b20f3264f0900100ba361d0082be0f00b9353264f2bf7e00b8341d0022b00c),
    .INIT_0E(256'h014808366410d02001490e1d0200900d0033013264f2d0010003801d0100300f),
    .INIT_0F(256'h0149080100209006000390207702203a02f80d050400900602f30c2076a3603f),
    .INIT_10(256'h0142062076a36046014308366480d0800142001d0400900d0149082265509006),
    .INIT_11(256'h014006226550900700b0020100209007001302207702204102f20e030bf09007),
    .INIT_12(256'h004300030bf207430140062076a20733014006360172074f0140061d08025000),
    .INIT_13(256'h00b43820113207510250002265520741037000010022075302f30f207702070f),
    .INIT_14(256'h01ba00207702075501b900050402070f0188402076a2072b001200208d52074d),
    .INIT_15(256'h02f935220082070b02f834207aa207130112012077c2070f03ac5c0100020715),
    .INIT_16(256'h022c51250003e05a032c7e366581900101c2d00d0800101902fa360900d25000),
    .INIT_17(256'h02f20f25000200c200ba363665c200dc00b9350d040200d400b8340900d25000),
    .INIT_18(256'h01b9000b215208c601884001300320600194020150a0d00100b438014400900d),
    .INIT_19(256'h00b93514300208e700b834142002090403ecab0d0100110101ba000b01401080),
    .INIT_1A(256'h02f30c0300701000001300143003606300b20f142001dc9300ba360d00820914),
    .INIT_1B(256'h014908141062f0020149083a67101000000390190012f00102f80d0110105001),
    .INIT_1C(256'h02f20e2d30a1d104014200123500311e01430810240001e00142002266d20bbb),
    .INIT_1D(256'h014006250001d112014006020103207c00b002090081d1060013032d2093207a),
    .INIT_1E(256'h02f30f14b062208700430014b06012020140060bb132201701400601a003207e),
    .INIT_1F(256'h00120009f1f0dd1000b40309e1e0100002500009d1d2208703700009c1c01206),
    .INIT_20(256'h03ac8913e000dd2001ba0013d001400001b90010cb00dd4001884010ba036085),
    .INIT_21(256'h02fa36206a22f23902f93501b000122102f83401a042f00201120113f0014000),
    .INIT_22(256'h00ba3609d070900200b935206582f03a00b83409c0701000022c8020658200be),
    .INIT_23(256'h01884009f07200ce019402206582f02400b40309e070100102f20f206580d004),
    .INIT_24(256'h00b8340b511208d503ecab0b410208cf01ba0001b01208d201b90001a73200e7),
    .INIT_25(256'h00130012d502093d00b20f10c402b02e00ba36036012093d00b9350b6122b02e),
    .INIT_26(256'h0149081bb002010500039019a01200c802f80d13f00200be02f30c12e60208c6),
    .INIT_27(256'h01420001b010300f01430801a7409001014200250002b04e0149083e696200be),
    .INIT_28(256'h0140062df070d00200b0022065c0900200130425000320b302f20e206a21d001),
    .INIT_29(256'h0043002dd072b40f0140062065c2b20f0140062de07208d50140062065c320ad),
    .INIT_2A(256'h0012ff2db07207aa0250002065c2077c0370002dc070100202f30f2065c2b80f),
    .INIT_2B(256'h02f20f0146c0100002f20e25000208d502f20d2da072011302f20c2065c22008),
    .INIT_2C(256'h00b0160b014208d50013000b2152200802500001300207aa037000015002077c),
    .INIT_2D(256'h02f1170d0080100102f016143002b80f020ccf142002b40f00b1170d0102b20f),
    .INIT_2E(256'h00b119011012071100b0180300720731001301143002079802f220142002f032),
    .INIT_2F(256'h02f221226bc2073f02f119141062074702f0183a6c0224b4020ccf190012070d),
    .INIT_30(256'h020ccf2d2092072f00b11b2d30a2073b00b01a1235025000001302102402070b),
    .INIT_31(256'h0013032d2092500002f2222d30a2070d02f11b060102074902f01a090082072b),
    .INIT_32(256'h02f01c14b0020751020ccf14a062073b00b11d250002074500b01c2d0082073b),
    .INIT_33(256'h00120014f002073102500014e002074d02f22314d002500002f11d14c002070d),
    .INIT_34(256'h01400614d082500003100014e082070d01f1ff14f0e2073f01d0ff250002072d),
    .INIT_35(256'h014100250000900101400614a082070d01400614b082074f01400614c0820735),
    .INIT_36(256'h01400e390002500001400e190e92070b01410039000206e4014006110b90300f),
    .INIT_37(256'h025000390000900200b224110072070d0100303e6e22073501400e190112072b),
    .INIT_38(256'h022ffd250001400e022ffd1100a1400e022ffd250001400e022ffd190f603008),
    .INIT_39(256'h022ffd2075f010c0022ffd206f625000022ffd206ec2070b022ffd00c00206e4),
    .INIT_3A(256'h022ffd2500001e00022ffd2075f01f00022ffd206f620904022ffd206ec01100),
    .INIT_3B(256'h022ffd14c06010a0022ffd141002091e022ffd14c0601c00022ffd0110001d01),
    .INIT_3C(256'h022ffd14c0601e00022ffd1410001f00022ffd14c0620904022ffd1410001100),
    .INIT_3D(256'h022ffd3a6f9010c0022ffd1d10a2091e022ffd2500001c00022ffd1410001d00),
    .INIT_3E(256'h022ffd01a0003f81022ffd250002091b022ffd1113020904022ffd1110701101),
    .INIT_3F(256'h022ffd3900005f00022ffd206d803c3f022ffd0900603d7c022ffd2076203e3c),
    .INIT_40(256'h022ffd367012091e022ffd1910105c00022ffd206ca05d03022ffd0110405e40),
    .INIT_41(256'h022ffd2075f20904022ffd206f601101022ffd00100010c0022ffd04a0025000),
    .INIT_42(256'h022ffd0110d03dfd022ffd2500003e7f022ffd366fc03fff022ffd192012091b),
    .INIT_43(256'h022ffd0115f05d00022ffd2275f05e80022ffd0112005f00022ffd2275f03cff),
    .INIT_44(256'h022ffd01131010c0022ffd2275f25000022ffd0113e2091e022ffd2275f05c00),
    .INIT_45(256'h022ffd0113003fff022ffd2275f2091b022ffd0113320904022ffd2275f01101),
    .INIT_46(256'h022ffd011322091e022ffd2275f03cff022ffd0113103dfe022ffd2275f03eff),
    .INIT_47(256'h022ffd0113420904022ffd2275f01101022ffd01133010c0022ffd2275f25000),
    .INIT_48(256'h022ffd0113603dfe022ffd2275f03eff022ffd0113503fff022ffd2275f2091b),
    .INIT_49(256'h022ffd0113805d01022ffd2275f05e00022ffd0113705f00022ffd2275f03cff),
    .INIT_4A(256'h022ffd0114101000022ffd2275f25000022ffd011392091e022ffd2275f05c00),
    .INIT_4B(256'h022ffd011430d040022ffd2275f0900f022ffd011422f01e022ffd2275f2f032),
    .INIT_4C(256'h022ffd011450d080022ffd2275f36171022ffd011440d020022ffd2275f36171),
    .INIT_4D(256'h022ffd0114736168022ffd2275f0d080022ffd011460900e022ffd2275f3616c),
    .INIT_4E(256'h022ffd0114936162022ffd2275f0d020022ffd0114836165022ffd2275f0d040),
    .INIT_4F(256'h022ffd0114b0d004022ffd2275f0900e022ffd0114a3615f022ffd2275f0d010),
    .INIT_50(256'h022ffd0114d2b04e022ffd2275f2f033022ffd0114c09016022ffd2275f32148),
    .INIT_51(256'h022ffd0114f22156022ffd2275f36155022ffd0114e1d00e022ffd2275f0300f),
    .INIT_52(256'h022ffd0115109006022ffd2275f36155022ffd011500d020022ffd2275f0900d),
    .INIT_53(256'h022ffd011531d053022ffd2275f22156022ffd011523614f022ffd2275f1d049),
    .INIT_54(256'h022ffd01155207b3022ffd2275f2070b022ffd011542074f022ffd2275f36155),
    .INIT_55(256'h022ffd011572070b022ffd2275f2073b022ffd0115622008022ffd2275f207aa),
    .INIT_56(256'h022ffd0115901000022ffd2275f208d5022ffd0115820113022ffd2275f208c6),
    .INIT_57(256'h022ffd207662b10e022ffd2275f22008022ffd0115a207aa022ffd2275f2077c),
    .INIT_58(256'h022ffd0d02001040022ffd0900d2b20e022ffd250002216f022ffd2d10601080),
    .INIT_59(256'h022ffd0d0102216f022ffd0900d01020022ffd250002b40e022ffd367622216f),
    .INIT_5A(256'h022ffd030602216f022ffd0900001010022ffd250002b80e022ffd36766208c6),
    .INIT_5B(256'h022ffd250002f01e022ffd0309f01008022ffd090002b80f022ffd25000208c6),
    .INIT_5C(256'h022ffd041002b20f022ffd2076d2b40f022ffd03160208c6022ffd00100221e8),
    .INIT_5D(256'h022ffd2070d19801022ffd2072f0982f022ffd207352f01e022ffd2d10001001),
    .INIT_5E(256'h022ffd2500020904022ffd2070b01102022ffd206e4010a0022ffd2076a0b237),
    .INIT_5F(256'h022ffd041002fc0c022ffd2076a03f07022ffd0319f20914022ffd00100208e7),
    .INIT_60(256'h022ffd2070d0bc0c022ffd2072f2ff0f022ffd2074f2fe0e022ffd2d1002fd0d),
    .INIT_61(256'h022ffd2076d01020022ffd327a60bf0f022ffd1d0010be0e022ffd0b0320bd0d),
    .INIT_62(256'h022ffd2074f0b001022ffd250002091e022ffd2070b20904022ffd206e401100),
    .INIT_63(256'h022ffd206e422193022ffd0100222017022ffd2070d36190022ffd2072f0d001),
    .INIT_64(256'h022ffd0319f0b016022ffd0010020941022ffd25000208f3022ffd2070b208db),
    .INIT_65(256'h022ffd250000b018022ffd2d1001f000022ffd041000b017022ffd2076a1d000),
    .INIT_66(256'h022ffd2d1030b01a022ffd0b1321f000022ffd207920b019022ffd010001f000),
    .INIT_67(256'h022ffd0b0320b01c022ffd2070d1f000022ffd2072f0b01b022ffd2074f1f000),
    .INIT_68(256'h022ffd206e4361af022ffd010401f000022ffd327a60b01d022ffd1d0011f000),
    .INIT_69(256'h022ffd206e40b03a022ffd0102032507022ffd250001d002022ffd2070b0b032),
    .INIT_6A(256'h022ffd1d0000b032022ffd2076d208d5022ffd250002f03a022ffd2070b11001),
    .INIT_6B(256'h022ffd2070d0b001022ffd2071122008022ffd20747324b4022ffd327b11d001),
    .INIT_6C(256'h022ffd2074f321e5022ffd227ae1d800022ffd2073b3092a022ffd250000d001),
    .INIT_6D(256'h022ffd206e52f035022ffd0bc020b017022ffd2070d2f034022ffd207450b016),
    .INIT_6E(256'h022ffd2074d2f03b022ffd207750b019022ffd207812f036022ffd2070b0b018),
    .INIT_6F(256'h022ffd206e52f03d022ffd0bc3a0b01b022ffd2070d2f03c022ffd2073b0b01a),
    .INIT_70(256'h022ffd207352f03f022ffd207430b01d022ffd250002f03e022ffd2070b0b01c),
    .INIT_71(256'h022ffd0bc0620941022ffd20717208f3022ffd20717208db022ffd2070d20921),
    .INIT_72(256'h022ffd0bc040b017022ffd206e51c010022ffd0bc050b134022ffd206e50b016),
    .INIT_73(256'h022ffd207510b136022ffd208180b018022ffd2070b1e010022ffd206e50b135),
    .INIT_74(256'h022ffd0d5041e010022ffd095020b13b022ffd2070d0b019022ffd2072d1e010),
    .INIT_75(256'h022ffd09c1c0b01b022ffd227ee1e010022ffd2082a0b13c022ffd3a7d70b01a),
    .INIT_76(256'h022ffd0bb020b13e022ffd09f1f0b01c022ffd09e1e1e010022ffd09d1d0b13d),
    .INIT_77(256'h022ffd13d001e010022ffd10cb00b13f022ffd14b060b01d022ffd14b061e010),
    .INIT_78(256'h022ffd2fe36321e5022ffd2ff3b1d800022ffd13f0019801022ffd13e00361f7),
    .INIT_79(256'h022ffd206e52f01f022ffd0bc3b01004022ffd2fc3420ae1022ffd2fd35221c4),
    .INIT_7A(256'h022ffd206e51d002022ffd0bc350b032022ffd206e52f013022ffd0bc360b002),
    .INIT_7B(256'h022ffd2072f0b032022ffd2070b207bb022ffd206e52070b022ffd0bc34321ee),
    .INIT_7C(256'h022ffd3a7f63252b022ffd0d5041d002022ffd2070d3252b022ffd2072d1d001),
    .INIT_7D(256'h022ffd0bd350b03a022ffd0bc3422008022ffd2280c2077c022ffd2082a01004),
    .INIT_7E(256'h022ffd01b001d000022ffd01a040b016022ffd0bf3b2f03a022ffd0be3611001),
    .INIT_7F(256'h022ffd206581f000022ffd09f070b018022ffd206581f000022ffd206a20b017),
    .INITP_00(256'ha73329e315aa3dd7ede220811bbeac5fab0537a82ab51610b312c2e5e7a41131),
    .INITP_01(256'h85a178fdaf29af2e163bb0a3f73c8a288b2fdf0c8cab454628ed65772be01da6),
    .INITP_02(256'hd61cb732e677ad4652e820cab6382880bf6867e4082b913f383226e5039b9185),
    .INITP_03(256'h1da3e7cafa8f15b8a52e121849001111091122c849b02300231ecb3d10bd8413),
    .INITP_04(256'ha0a214378da3efd12299a3811f7515150e27397b0fb434db54c26231dd820bb6),
    .INITP_05(256'h5e6a4178af31077e4767702321ae78f7ce61d3ee3046c5d00c9abc860418bcc3),
    .INITP_06(256'hcf0c0f03aa9622ad13872a02ade497ae9ef0e575ccc3a60591e9e7f4e080a230),
    .INITP_07(256'hc86fc8616ff8fa774d75f7f95df752e74bfe535ff9e7fc767de0f347fd55fd7c),
    .INITP_08(256'h4ddc4851c15cd4524343d0dcd35140d8775a595cd265c2c2e56defe3e1de625c),
    .INITP_09(256'h7543f45a7459eed8ec5ff8cb6540794065c07dd17451ddd8d7d65a5c49524543),
    .INITP_0A(256'h6443fb5277cdea42e5d9665ff6dae94c62c87e4afc4cfb45f44ce7c66b527053),
    .INITP_0B(256'hdbf3cd71f651e0f64f53ca635979c979617f41f9e74fedc66cd7f3d7fbc6f4eb),
    .INITP_0C(256'h7ada54e06cd3696861644eead779ff42fe68c2d8e1fdc6eb6a604c63c74575f4),
    .INITP_0D(256'hf864d955f8e87851fff9deee61ccdfebdb507febc47f6d4c61f1fb59fec971da),
    .INITP_0E(256'h504f627058d27ae954f4d1e16a5255deebca46f17e70e570fbd05dcec368ebd7),
    .INITP_0F(256'hc057c0cfdafef35a4ee168dee0e757555ade74f4ee6a76e8f776e1d6cf747ad5),
